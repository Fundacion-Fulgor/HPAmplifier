* Extracted by KLayout with SG13G2 LVS runset on : 23/01/2026 16:17

.SUBCKT OTA_Telescopic_CMFB VSS VINP VINN CMFB VREF VDD IBIAS
M$1 CMFB CMFB VSS VSS sg13_lv_nmos L=0.2u W=29.97u AS=6.1938p AD=5.6943p
+ PS=37.02u PD=33.39u
M$10 VSS \$5 \$5 VSS sg13_lv_nmos L=0.2u W=29.97u AS=5.6943p AD=6.1938p
+ PS=33.39u PD=37.02u
M$19 \$5 VREF \$42 VDD sg13_lv_pmos L=0.35u W=35.98u AS=7.2217p AD=6.8362p
+ PS=49.79u PD=46.62u
M$33 \$5 VREF \$64 VDD sg13_lv_pmos L=0.35u W=35.98u AS=6.8362p AD=7.2217p
+ PS=46.62u PD=49.79u
M$47 CMFB VINP \$42 VDD sg13_lv_pmos L=0.35u W=35.98u AS=7.2217p AD=6.8362p
+ PS=49.79u PD=46.62u
M$61 CMFB VINN \$64 VDD sg13_lv_pmos L=0.35u W=35.98u AS=6.8362p AD=7.2217p
+ PS=46.62u PD=49.79u
M$75 VDD IBIAS \$42 VDD sg13_lv_pmos L=0.7u W=144u AS=28.26p AD=27.36p
+ PS=206.52u PD=198.72u
M$99 VDD IBIAS \$64 VDD sg13_lv_pmos L=0.7u W=144u AS=27.36p AD=28.26p
+ PS=198.72u PD=206.52u
M$419 VDD IBIAS IBIAS VDD sg13_lv_pmos L=0.7u W=48u AS=9.27p AD=9.27p PS=67.54u
+ PD=67.54u
.ENDS OTA_Telescopic_CMFB
