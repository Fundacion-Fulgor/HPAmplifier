** sch_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_TOP_TB_OL.sch
**.subckt OTA_Telescopic_TOP_TB_OL
V7 net1 GND 1.25
C1 Vout1 GND 500f m=1
C2 Vout2 GND 500f m=1
x1 VDD GND net3 net1 net4 Vout2 Vout1 net1 net2 net1 VREF net5 net5 OTA_Telescopic_TOP
V6 VDD GND 1.8
R3 net3 net4 10G m=1
R4 net2 net1 10G m=1
V1 net4 net1 0 AC 1
V2 VREF GND dc 0.9 pwl(0 0.8 1u 0.8 1.01u 0.9 0.15m 0.9 0.15m 0)
**** begin user architecture code

** opencircuitdesign pdks install
.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ
.lib cornerCAP.lib cap_typ
.temp 65



.control
save all
 set color0 = white

* AC simulation
ac dec 1k 1 1T
let Av = db((v(Vout2)-v(Vout1)))
meas ac Ao FIND Av WHEN frequency=10
let ABW = Ao-3
meas ac BW WHEN Av=ABW
meas ac UGBW WHEN Av=0
let phase_vec = 180/pi*cph(v(Vout2)-v(Vout1))

* Phase margin (PM)
meas ac phase FIND phase_vec WHEN frequency=UGBW
let PM = phase+180
print PM

* Gain margin (GM)
meas ac freq180 FIND frequency WHEN phase_vec=-180
meas ac gain FIND Av WHEN frequency=freq180
let GM = 0-gain

*BW in 7 dB
meas ac UGBW7dB WHEN Av=7
meas ac UGBW4dB WHEN Av=4

print GM
plot Av
plot phase_vec

plot db(v(x1.Vo1)-v(x1.Vo2))

write AC_OL.raw

wrdata AvOL_ Av
wrdata PhaseOL_ phase_vec


*DC simulation

op
let vout_dc = v(Vout1)
print vout_dc
write OTA_Telescopic_TOP_TB_OL.raw


reset
noise v(Vout1) V6 dec 100 1 0.5e9 1
setplot noise1
*plot onoise_spectrum
setplot noise2
print onoise_total

.endc


**** end user architecture code
**.ends

* expanding   symbol:  OTA_Telescopic_TOP.sym # of pins=13
** sym_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_TOP.sym
** sch_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_TOP.sch
.subckt OTA_Telescopic_TOP VDD VSS VPout VP VPin VOUTN VOUTP VNin VNout VN VREF CMFBin CMFBout
*.ipin VP
*.ipin VN
*.opin VOUTP
*.opin VOUTN
*.ipin VPin
*.ipin VNin
*.opin VPout
*.opin VNout
*.iopin VDD
*.iopin VSS
*.iopin VREF
*.ipin CMFBin
*.opin CMFBout
x1 VDD CMFBin VOUTN VOUTP VPin VNin VSS net2 OTA_Telescopic_core
x2 VDD VREF VOUTN VOUTP net1 CMFBout VSS OTA_Telescopic_CMFB
XM3 net2 vbp VDD VDD sg13_lv_pmos w=12u l=2.5u ng=2 m=1
XM2 net1 vbn VSS VSS sg13_lv_nmos w=12.5u l=6.5u ng=2 m=1
XR3 VN VNout VSS rppd w=0.6e-6 l=6.73e-6 m=1 b=0
XR4 VPout VP VSS rppd w=0.6e-6 l=6.73e-6 m=1 b=0
XR5 VOUTP VPout VSS rppd w=0.6e-6 l=15.4e-6 m=1 b=0
XR2 VOUTN VNout VSS rppd w=0.6e-6 l=15.4e-6 m=1 b=0
x3 VDD vbp vbn VSS OTA_Telescopic_currentRef
.ends


* expanding   symbol:  OTA_Telescopic_core.sym # of pins=8
** sym_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_core.sym
** sch_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_core.sch
.subckt OTA_Telescopic_core VDD CMFB VOUTP VOUTN VINP VINN VSS IB
*.iopin VDD
*.iopin VSS
*.ipin VINP
*.ipin VINN
*.opin VOUTN
*.opin VOUTP
*.ipin CMFB
*.iopin IB
V2 VB2 VSS 1.5
V3 VB3 VSS 0.7
V4 VB4 VSS 0.49409
V1 VB5 VSS 1.15
* noconn VB2
* noconn VB3
* noconn VB4
* noconn VB5
V5 VB VSS 0.90204
* noconn VB
XM15 VB55 VB55 VDD VDD sg13_lv_pmos w=1.4u l=0.35u ng=1 m=8
XM17 VB33 VB33 VDD VDD sg13_lv_pmos w=2.05u l=0.35u ng=1 m=1
XM18 VB22 VB33 VDD VDD sg13_lv_pmos w=2.05u l=0.35u ng=1 m=1
XM9 VOUTP Vo1 VDD VDD sg13_lv_pmos w=1.37u l=0.35u ng=1 m=200
XM7 Vx1 VB55 VDD VDD sg13_lv_pmos w=7u l=0.7u ng=1 m=30
XM5 Vo1 VB33 Vx1 VDD sg13_lv_pmos w=4.05u l=0.5u ng=1 m=30
XM8 Vx2 VB55 VDD VDD sg13_lv_pmos w=7u l=0.7u ng=1 m=30
XM6 Vo2 VB33 Vx2 VDD sg13_lv_pmos w=4.05u l=0.5u ng=1 m=30
XM10 VOUTN Vo2 VDD VDD sg13_lv_pmos w=1.37u l=0.35u ng=1 m=200
XM13 IB IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM14 VB55 IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM16 VB33 IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM19 VB22 VB22 VSS VSS sg13_lv_nmos w=0.5u l=0.8u ng=1 m=1
XM11 VOUTP IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=55
XM0 P CMFB VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=34
XM3 Vo1 VB22 Vy1 VSS sg13_lv_nmos w=1.9u l=0.16u ng=1 m=30
XM1 Vy1 VINP P VSS sg13_lv_nmos w=1.1u l=0.15u ng=1 m=30
XM4 Vo2 VB22 Vy2 VSS sg13_lv_nmos w=1.9u l=0.16u ng=1 m=30
XM2 Vy2 VINN P VSS sg13_lv_nmos w=1.1u l=0.15u ng=1 m=30
XM12 VOUTN IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=55
XR3 VOUTP net1 VSS rppd w=1.3e-6 l=0.55e-6 m=1 b=0
XR1 net2 VOUTN VSS rppd w=1.3e-6 l=0.55e-6 m=1 b=0
XC3 Vo2 net2 cap_cmim w=21e-6 l=21e-6 m=1
XC1 Vo1 net1 cap_cmim w=21e-6 l=21e-6 m=1
.ends


* expanding   symbol:  OTA_Telescopic_CMFB.sym # of pins=7
** sym_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_CMFB.sym
** sch_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_CMFB.sch
.subckt OTA_Telescopic_CMFB VDD VREF VINN VINP IBIAS CMFB VSS
*.iopin VDD
*.iopin VSS
*.opin CMFB
*.ipin VREF
*.iopin IBIAS
*.ipin VINP
*.ipin VINN
XM0 IBIAS IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=8
XM1 V1 IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=24
XM2 V2 IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=24
XM3 CMFB VINP V1 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM4 net1 VREF V1 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM5 net1 VREF V2 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM6 CMFB VINN V2 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM7 net1 net1 VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=6
XM8 CMFB CMFB VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=6
.ends


* expanding   symbol:  OTA_Telescopic_currentRef.sym # of pins=4
** sym_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_currentRef.sym
** sch_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/HPAmplifier/OTA_Telescopic/OTA_Telescopic_currentRef.sch
.subckt OTA_Telescopic_currentRef VDD OUT_P OUT_N VSS
*.iopin VDD
*.iopin VSS
*.opin OUT_P
*.opin OUT_N
XM3 OUT_P OUT_P VDD VDD sg13_lv_pmos w=12u l=2.5u ng=2 m=1
XM2 OUT_P OUT_N net1 VSS sg13_lv_nmos w=12u l=6.4u ng=2 m=8
XM4 OUT_N OUT_P VDD VDD sg13_lv_pmos w=12u l=2.5u ng=2 m=1
XM1 OUT_N OUT_N VSS VSS sg13_lv_nmos w=12u l=6.4u ng=2 m=1
XM5 OUT_P OUT_P OUT_N VSS sg13_lv_nmos w=2u l=1u ng=1 m=1
XR2 VSS net1 VSS rppd w=1e-6 l=13.5e-6 m=1 b=0
.ends

.GLOBAL GND
.end
