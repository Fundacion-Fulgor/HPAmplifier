** sch_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/OTA_Telescopic_TOP_TB_CL.sch
**.subckt OTA_Telescopic_TOP_TB_CL
V7 net1 GND 1.25
V5 VP net1 0 SIN(0 0.0558 100000000) AC 0.5
V1 VDD GND 1.62
V2 VREF GND dc 0.9
C1 Vout1 GND 500f m=1
C2 Vout2 GND 500f m=1
V3 net1 VN 0 SIN(0 0.0558 100000000) AC 0.5
x1 VDD GND net2 VP net2 Vout2 Vout1 net3 net3 VN VREF net4 net4 OTA_Telescopic_TOP
**** begin user architecture code

** opencircuitdesign pdks install
.lib cornerMOSlv.lib mos_ss
.lib cornerRES.lib res_typ
.temp 125



.control
save all
 set color0 = white

* AC simulation
ac dec 1000 1 1T
let Av = db(v(Vout1)-v(Vout2))
meas ac Ao FIND Av WHEN frequency=10
let ABW = Ao-3
meas ac BW WHEN Av=ABW
meas ac UGBW WHEN Av=0
let phase_vec = 180/pi*cph(v(Vout1)-v(Vout2))

* Phase margin (PM)
meas ac phase FIND phase_vec WHEN frequency=UGBW
let PM = phase+180
print PM

* Gain margin (GM)
meas ac freq180 FIND frequency WHEN phase_vec=-180
meas ac gain FIND Av WHEN frequency=freq180
let GM = 0-gain

print GM
plot Av
plot phase_vec

write AC_OL.raw
wrdata AvCL_ Av

*DC simulation

op
let vout_dc = v(Vout1)
print vout_dc
write OTA_Telescopic_TB2_CL.raw

.endc


**** end user architecture code
**.ends

* expanding   symbol:  OTA_Telescopic_TOP.sym # of pins=13
** sym_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/OTA_Telescopic_TOP.sym
** sch_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/OTA_Telescopic_TOP.sch
.subckt OTA_Telescopic_TOP VDD VSS VPout VP VPin VOUTN VOUTP VNin VNout VN VREF CMFBin CMFBout
*.ipin VP
*.ipin VN
*.opin VOUTP
*.opin VOUTN
*.ipin VPin
*.ipin VNin
*.opin VPout
*.opin VNout
*.iopin VDD
*.iopin VSS
*.iopin VREF
*.ipin CMFBin
*.opin CMFBout
R5 VPout VP 3k m=1
R6 VNout VN 3k m=1
x1 VDD CMFBin VOUTN VOUTP VPin VNin VSS net2 OTA_Telescopic_core_v2
x2 VDD VREF VOUTN VOUTP net1 CMFBout VSS OTA_Telescopic_CMFB2
R1 VOUTN VNout 6.72k m=1
R2 VOUTP VPout 6.72k m=1
XM3 net2 vbp VDD VDD sg13_lv_pmos w=22u l=2u ng=4 m=1
XM2 net1 vbn VSS VSS sg13_lv_nmos w=9.86u l=9.86u ng=1 m=1
x3 VDD vbp vbn VSS currentRef
.ends


* expanding   symbol:  OTA_Telescopic_core_v2.sym # of pins=8
** sym_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/OTA_Telescopic_core_v2.sym
** sch_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/OTA_Telescopic_core_v2.sch
.subckt OTA_Telescopic_core_v2 VDD CMFB VOUTP VOUTN VINP VINN VSS IB
*.iopin VDD
*.iopin VSS
*.ipin VINP
*.ipin VINN
*.opin VOUTN
*.opin VOUTP
*.ipin CMFB
*.iopin IB
V2 VB2 VSS 1.5
V3 VB3 VSS 0.7
V4 VB4 VSS 0.49409
V1 VB5 VSS 1.12
* noconn VB2
* noconn VB3
* noconn VB4
* noconn VB5
V5 VB VSS 0.90204
* noconn VB
R1 net1 VOUTP 190 m=1
R2 VOUTN net2 190 m=1
C1 Vo1 net1 0.7p m=1
C2 Vo2 net2 0.7p m=1
XM15 VB55 VB55 VDD VDD sg13_lv_pmos w=1.45u l=0.35u ng=1 m=6
XM17 VB33 VB33 VDD VDD sg13_lv_pmos w=2.05u l=0.35u ng=1 m=1
XM18 VB22 VB33 VDD VDD sg13_lv_pmos w=2.05u l=0.35u ng=1 m=1
XM9 VOUTP Vo1 VDD VDD sg13_lv_pmos w=2u l=0.35u ng=1 m=250
XM7 Vx1 VB55 VDD VDD sg13_lv_pmos w=6.85u l=0.7u ng=1 m=30
XM5 Vo1 VB33 Vx1 VDD sg13_lv_pmos w=4.3u l=0.5u ng=1 m=30
XM8 Vx2 VB55 VDD VDD sg13_lv_pmos w=6.85u l=0.7u ng=1 m=30
XM6 Vo2 VB33 Vx2 VDD sg13_lv_pmos w=4.3u l=0.5u ng=1 m=30
XM10 VOUTN Vo2 VDD VDD sg13_lv_pmos w=2u l=0.35u ng=1 m=250
XM13 IB IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM14 VB55 IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM16 VB33 IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM19 VB22 VB22 VSS VSS sg13_lv_nmos w=0.5u l=0.8u ng=1 m=1
XM11 VOUTP IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=55
Xq P CMFB VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=43
XM3 Vo1 VB22 Vy1 VSS sg13_lv_nmos w=1.9u l=0.16u ng=1 m=30
XM1 Vy1 VINP P VSS sg13_lv_nmos w=1.1u l=0.15u ng=1 m=30
XM4 Vo2 VB22 Vy2 VSS sg13_lv_nmos w=1.9u l=0.16u ng=1 m=30
XM2 Vy2 VINN P VSS sg13_lv_nmos w=1.1u l=0.15u ng=1 m=30
XM12 VOUTN IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=55
.ends


* expanding   symbol:  OTA_Telescopic_CMFB2.sym # of pins=7
** sym_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/OTA_Telescopic_CMFB2.sym
** sch_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/OTA_Telescopic_CMFB2.sch
.subckt OTA_Telescopic_CMFB2 VDD VREF VINN VINP IBIAS CMFB VSS
*.iopin VDD
*.iopin VSS
*.opin CMFB
*.ipin VREF
*.iopin IBIAS
*.ipin VINP
*.ipin VINN
XM0 IBIAS IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=8
XM1 V1 IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=24
XM2 V2 IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=24
XM3 CMFB VINP V1 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=24
XM4 net1 VREF V1 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=24
XM5 net1 VREF V2 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=24
XM6 CMFB VINN V2 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=24
XM7 net1 net1 VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=8
XM8 CMFB CMFB VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=8
.ends


* expanding   symbol:  currentRef.sym # of pins=4
** sym_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/currentRef.sym
** sch_path: /foss/designs/HPAmplifier/Differential_OTA_Telescopic_IHP/currentRef.sch
.subckt currentRef VDD OUT_P OUT_N VSS
*.iopin VDD
*.iopin VSS
*.opin OUT_P
*.opin OUT_N
XM3 OUT_P OUT_P VDD VDD sg13_lv_pmos w=22u l=2u ng=4 m=1
XM2 OUT_P OUT_N net1 net1 sg13_lv_nmos w=9.86u l=9.86u ng=1 m=15
XM4 OUT_N OUT_P VDD VDD sg13_lv_pmos w=22u l=2u ng=4 m=1
XM1 OUT_N OUT_N VSS VSS sg13_lv_nmos w=9.86u l=9.86u ng=1 m=1
XM5 OUT_P OUT_P OUT_N VSS sg13_lv_nmos w=1u l=1u ng=1 m=1
XR2 VSS net1 sub! rppd w=0.6e-6 l=14e-6 m=1 b=0
.ends

.GLOBAL GND
.end
